////////////////////////////////////////////////////////////////////////////////
// Filename    : ahb_interconnect_compare.sv
// Description : 
//
// Author      : Phu Vuong
// History     : Mar 26, 2024 : Initial     
//
////////////////////////////////////////////////////////////////////////////////
module ahb_interconnect_compare_1bit (
    output logic    ol,
    output logic    oe,
    input           fl, //flag larger
    input           fe, //flag equal
    input           a,
    input           b
);
    ////////////////////////////////////////////////////////////////////////////
    //design description
    ////////////////////////////////////////////////////////////////////////////
    assign ol = fl | a | ~b;
    assign oe = a ~^ b;
endmodule